// ============================================================================
//        __
//   \\__/ o\    (C) 2009-2024  Robert Finch, Waterloo
//    \  __ /    All rights reserved.
//     \/_//     robfinch<remove>@finitron.ca
//       ||
//
// CALL NEAR Indirect
//
// BSD 3-Clause License
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this
//    list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
//
// 3. Neither the name of the copyright holder nor the names of its
//    contributors may be used to endorse or promote products derived from
//    this software without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
// FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
// DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
// OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// ============================================================================

rf80386_pkg::CALL_IN:
	begin
		if (StkAddrSize==8'd32) begin
			if (OperandSize32)
				esp <= esp - 4'd4;
			else
				esp <= esp - 4'd2;
		end
		else begin
			if (OperandSize32)
				esp[15:0] <= esp - 4'd4;
			else
				esp[15:0] <= esp - 4'd2;
		end
		tGoto(rf80386_pkg::CALL_IN1);
	end
rf80386_pkg::CALL_IN1:
	begin
		ad <= sssp;
		dat <= eip;
		sel <= OperandSize32 ? 16'h000F: 16'h0003;
		tGosub(rf80386_pkg::STORE,rf80386_pkg::CALL_IN2);
	end
rf80386_pkg::CALL_IN2:
	begin
		if (OperandSize32) begin
			ea <= cs_base + b;
			if (mod==2'b11) begin
				eip <= b;
				tGoto(rf80386_pkg::IFETCH);
			end
			else 
				tGoto(rf80386_pkg::CALL_IN3);
		end
		else begin
			ea <= cs_base + b[15:0];
			if (mod==2'b11) begin
				eip <= b[15:0];
				tGoto(rf80386_pkg::IFETCH);
			end
			else 
				tGoto(rf80386_pkg::CALL_IN3);
		end
	end
rf80386_pkg::CALL_IN3:
	begin
		ad <= ea;
		if (OperandSize32)
			sel <= 16'h000F;
		else
			sel <= 16'h0003;
		tGosub(rf80386_pkg::LOAD,rf80386_pkg::CALL_IN4);
	end
rf80386_pkg::CALL_IN4:
	begin
		if (OperandSize32)
			b[31:0] <= dat[31:0];
		else
			b[15:0] <= dat[15:0];
		tGoto(rf80386_pkg::CALL_IN5);
	end
rf80386_pkg::CALL_IN5:
	begin
		if (OperandSize32)
			eip <= b;
		else
			eip <= b[15:0];
		tGoto(rf80386_pkg::IFETCH);
	end
