// ============================================================================
//        __
//   \\__/ o\    (C) 2009-2024  Robert Finch, Waterloo
//    \  __ /    All rights reserved.
//     \/_//     robfinch<remove>@finitron.ca
//       ||
//
//  BRANCH.v
//  Jcc disp8
//  - conditional branches
//  - fetch an 8 bit displacement and add into IP
//
// BSD 3-Clause License
// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this
//    list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright notice,
//    this list of conditions and the following disclaimer in the documentation
//    and/or other materials provided with the distribution.
//
// 3. Neither the name of the copyright holder nor the names of its
//    contributors may be used to endorse or promote products derived from
//    this software without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE
// FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
// DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER
// CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY,
// OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE
// OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// ============================================================================

// Fetch branch displacement if taking branch, otherwise skip

rf80386_pkg::BRANCH1:
	if (take_br) begin
		if (jccl) begin
			if (cs_desc.db) begin
				disp32 <= bundle[31:0];
				eip <= eip + 4'd4;
			end
			else begin
				disp32 <= {{16{bundle[15]}},bundle[15:0]};
				eip <= eip + 4'd2;
			end
		end
		else begin
			disp32 <= {{24{bundle[7]}},bundle[7:0]};
			eip <= eip + 4'd1;
		end
		tGoto(rf80386_pkg::BRANCH2);
	end
	else begin
		if (jccl) begin
			if (cs_desc.db)
				eip <= eip + 4'd4;
			else
				eip <= eip + 4'd2;
		end
		else
			eip <= eip + 4'd1;
		tGoto(rf80386_pkg::IFETCH);
	end
BRANCH2:
	begin
		eip <= eip + disp32;
		tGoto(rf80386_pkg::IFETCH);
	end
